library verilog;
use verilog.vl_types.all;
entity ELEVADOR_vlg_vec_tst is
end ELEVADOR_vlg_vec_tst;
